module yAdder1(z, cout, a, b, cin); 
	output z, cout; 
	input a, b, cin; 
	xor left_xor(tmp, a, b); 
	xor right_xor(z, cin, tmp); 
	and left_and(outL, a, b); 
	and right_and(outR, tmp, cin); 
	or my_or(cout, outR, outL); 
endmodule 
